LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MBR IS
	PORT(
		MBR_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		MBR_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		MEM_IN : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		MEM_OUT : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		R,W : IN STD_LOGIC
	);
END MBR;

ARCHITECTURE BEHAVI OF MBR IS
SIGNAL MBR_REG : STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
BEGIN
	PROCESS(R, W)
	BEGIN
		IF R = '1' THEN
			MBR_REG <= MEM_OUT; 
		ELSIF W = '1' THEN
			MBR_REG <= MBR_IN;
		END IF;
		MBR_OUT <= MBR_REG;
		MEM_IN <= MBR_REG;
	END PROCESS;
END;