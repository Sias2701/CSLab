LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MAR IS
	PORT(
		MAR_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		PEND : IN STD_LOGIC;
		MAR_OUT : BUFFER STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END MAR;

ARCHITECTURE BEHAVI OF MAR IS
SIGNAL MAR_REG : STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
	PROCESS(PEND)
	BEGIN
		IF PEND = '1' THEN
			MAR_REG <= MAR_IN;
		END IF;
		MAR_OUT <= MAR_REG;
	END PROCESS;
END BEHAVI;