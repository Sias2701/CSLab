LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY PC IS
	PORT(
		PC_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		PC_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		RST, PEND, INC: IN STD_LOGIC
	);
END PC;

ARCHITECTURE BEHAVI OF PC IS
SIGNAL PROGRAM_COUNTER_REG : STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
	PROCESS(RST)
	BEGIN
		IF RST = '1' THEN
			IF RISING_EDGE(PEND) THEN
				IF INC = '1' THEN
					PROGRAM_COUNTER_REG <= "00000001" + PROGRAM_COUNTER_REG;
				ELSE
					PROGRAM_COUNTER_REG <= PC_IN;
				END IF;
			END IF;
			PC_OUT <= PROGRAM_COUNTER_REG;
		ELSE
			PROGRAM_COUNTER_REG <= "00000000";
		END IF;
	END PROCESS;
END BEHAVI;