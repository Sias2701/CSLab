-- 正弦波发生器
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY SineGenerator IS
	PORT(
		CLK : IN STD_LOGIC;
		DOUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END ENTITY SineGenerator;
ARCHITECTURE DACC OF SineGenerator IS
	COMPONENT data_rom IS 
	PORT(address  : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
		  clock  : IN STD_LOGIC ;
		  q        : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)	);
	END COMPONENT;

	SIGNAL Q1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
BEGIN
	PROCESS(CLK)
	BEGIN
	IF CLK'EVENT AND CLK = '1' THEN Q1<=Q1+1;
	END IF;
	END PROCESS;
u1 : data_rom PORT MAP(address=>Q1, q => DOUT,clock=>CLK);
END; 

