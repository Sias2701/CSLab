-- HalfAdder.vhd
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY HalfAdder IS
	PORT(a, b : IN STD_LOGIC; s, c : OUT STD_LOGIC);
END ENTITY HalfAdder;
ARCHITECTURE one OF HalfAdder IS
BEGIN
	s <= a XOR b;
	c <= a AND b;
END ARCHITECTURE one;
