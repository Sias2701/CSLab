LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY CAR IS
	PORT(
		OPCODE : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		BADDR : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		CU_LOOPBACK : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		CADDR : BUFFER STD_LOGIC_VECTOR(7 DOWNTO 0);
		CLK, RST : IN STD_LOGIC
	);
END CAR;

ARCHITECTURE BEHAVI OF CAR IS
BEGIN
	PROCESS(RST)
	BEGIN
	IF RST = '1' THEN
		IF RISING_EDGE(CLK) THEN
			IF CU_LOOPBACK = "1000" THEN
				CADDR <= "00000001" + CADDR;
			ELSIF CU_LOOPBACK = "0100" THEN
				CADDR <= OPCODE + CADDR;
			ELSIF CU_LOOPBACK = "0010" THEN
				CADDR <= BADDR;
			END IF;
		END IF;
	ELSE
		CADDR <= "00000000";
	END IF;
	END PROCESS;
END BEHAVI;