LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY CONTROL_UNIT IS
	PORT(
		CONTROL_WORD : IN STD_LOGIC_VECTOR(41 DOWNTO 0);
		CONTROL_BUS : OUT STD_LOGIC_VECTOR(21 DOWNTO 0);
		LOOP_BACK : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		ALU_MODE : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		BADDR : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		ACC_ZF : IN STD_LOGIC
	);
END CONTROL_UNIT;

ARCHITECTURE BEHAVI OF CONTROL_UNIT IS
BEGIN
	ALU_MODE <= CONTROL_WORD(40 DOWNTO 37);
	LOOP_BACK <= CONTROL_WORD(33 DOWNTO 30) WHEN CONTROL_WORD(34) = '0' ELSE
					 "0010" WHEN (CONTROL_WORD(35) = '1' AND ACC_ZF = '0') OR (CONTROL_WORD(36) = '1' AND ACC_ZF = '1') ELSE
					 "1000";
	CONTROL_BUS <= CONTROL_WORD(29 DOWNTO 8);
	BADDR <= CONTROL_WORD(7 DOWNTO 0);
END BEHAVI;