LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ALU IS
	PORT(
		ALU_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		ACC_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		RESULT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		PEND : IN STD_LOGIC;
		MODE : IN STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END ALU;

ARCHITECTURE BEHAVI OF ALU IS
SIGNAL ALU_BUF : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL MUL_BUF : STD_LOGIC_VECTOR(15 DOWNTO 0);
BEGIN
	PROCESS(ACC_IN, MODE, ALU_IN)
	BEGIN
		IF PEND = '1' THEN
			ALU_BUF <= ALU_IN;
		END IF;
		IF MODE = "0001" THEN
			RESULT <= ACC_IN + ALU_BUF;
		ELSIF MODE = "0010" THEN
			RESULT <= ACC_IN - ALU_BUF;
		ELSIF MODE = "0011" THEN
			MUL_BUF <= ACC_IN * ALU_BUF;
			RESULT <= MUL_BUF(7 DOWNTO 0);
		ELSIF MODE = "0100" THEN
			RESULT <= ACC_IN AND ALU_BUF;
		ELSIF MODE = "0101" THEN
			RESULT <= ACC_IN OR ALU_BUF;
		ELSIF MODE = "0110" THEN
			RESULT <= NOT ACC_IN;
		ELSIF MODE = "0111" THEN
			RESULT <= ACC_IN XOR ALU_BUF;
		ELSIF MODE = "1000" THEN
			RESULT <= ACC_IN(6 DOWNTO 0) & '0';
		ELSIF MODE = "1001" THEN
			RESULT <= '0' & ACC_IN(7 DOWNTO 1);
		ELSIF MODE = "1110" THEN
			RESULT <= ACC_IN + "00000001";
		ELSIF MODE = "1111" THEN
			RESULT <= ACC_IN - "00000001";
		ELSE
			RESULT <= ACC_IN;
		END IF;
	END PROCESS;
END BEHAVI;